module unsigned_to_20b_signed(
	input [LENGTH-1:0] in,
	output [19:0] out
)

	parameter LENGTH = 4;
	

endmodule