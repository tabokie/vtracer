module ray_tracer_ceiling(
	input [27:0] init,
	input [27:0] dir,
	input object_in, // 10-10-10-10(bound)-10(position)-2(axis) = 52
	output [9:0] t_out
);

endmodule
