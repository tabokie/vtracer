module ray_tracer_sphere(
	input sphere;
	input 
)

endmodule