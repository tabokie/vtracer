module div(
	input [LENGTH-1:0] in_0,
	input [LENGTH-1:0] in_1,
	output [LENGTH-1:0] out
);

	

endmodule